module datapath(input [31:0] x1, x2, x3, x4, 
        input rst, clk, init, start , write_reg,
        output reg [15:0] max_index,
        output reg done);
    
endmodule