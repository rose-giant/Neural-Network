`include "PU.v"

module PU_TB();

    reg [31:0] x1, x2, x3, x4, w1, w2, w3, w4;
    wire [31:0] result; 
    
    PU PU_instance(x1, x2, x3, x4, w1, w2, w3, w4, result);

    initial begin
        $dumpfile("PU_TB.vcd");
        $dumpvars(0, PU_TB);

        #10;
        x1 = 32'b11111111000001010100100010000;
        x2 = 32'b00110000110000000110000100010;
        x3 = 32'b11111111000001010100100010000;
        x4 = 32'b00110000110000000110000100010;

        w1 = 32'b11111111000001010100100010000;
        w2 = 32'b00110000110000000110000100010;
        w3 = 32'b11111111000001010100100010000;
        w4 = 32'b00110000110000000110000100010;

        
        x1 = 32'b11111111000001010100100010000;
        x2 = 32'b00110000110000000110000100010;
        x3 = 32'b11111111000001010100100010000;
        x4 = 32'b00110000110000000110000100010;

        w1 = 32'b00110000110000000110000100010;
        w2 = 32'b11111111000001010100100010000;
        w3 = 32'b11111111000001010100100010000;
        w4 = 32'b00110000110000000110000100010;

        #10;
        x1 = 32'b11111111000001010100100010000;
        x2 = 32'b00110000110000000110000100010;
        x3 = 32'b00110000110000000110000100010;
        x4 = 32'b11111111000001010100100010000;

        w1 = 32'b11111111000001010100100010000;
        w2 = 32'b00110000110000000110000100010;
        w3 = 32'b11111111000001010100100010000;
        w4 = 32'b00110000110000000110000100010;
    end

endmodule